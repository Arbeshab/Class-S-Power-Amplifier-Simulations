.subckt CSGP_0805_885012007066_3R3nF 1 2
Rser 1 3 0.0386718470366
Lser 2 4 4.52637868E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends CSGP_0805_885012007066_3R3nF