.subckt CSGP_1210_885012109011_47uF 1 2
Rser 1 3 0.00225907860771
Lser 2 4 0.0000000009
C1 3 4 0.000047
Rpar 3 4 1000000
.ends CSGP_1210_885012109011_47uF