.subckt CSGP_0805_885012007041_1R5nF 1 2
Rser 1 3 0.0403337213614
Lser 2 4 2.897145E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends CSGP_0805_885012007041_1R5nF