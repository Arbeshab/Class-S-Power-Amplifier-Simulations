.subckt ASLI_865080353015_470uF 1 2
Rser 1 3 0.133
Lser 2 4 2.09657010043051E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends ASLI_865080353015_470uF