.subckt ASLI_865080542005_15uF 1 2
Rser 1 3 0.89
Lser 2 4 1.787806959E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends ASLI_865080542005_15uF