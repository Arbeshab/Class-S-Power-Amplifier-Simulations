.subckt CBF_1806_74279246_1000ohm 1 2
Rp 1 2 1045
Cp 1 2 1.241p
Rs 1 N3 0.056
L1 N3 2 0.108u
.ends CBF_1806_74279246_1000ohm