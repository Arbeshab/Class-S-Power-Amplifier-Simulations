.subckt 865080653016_100uF 1 2
Rser 1 3 0.197
Lser 2 4 4.80864427233527E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080653016_100uF