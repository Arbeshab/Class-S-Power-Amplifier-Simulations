.subckt CSGP_0805_885012207097_68nF 1 2
Rser 1 3 0.0207501013107
Lser 2 4 0.00000000038
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends CSGP_0805_885012207097_68nF