.subckt CSGP_0805_885012007043_3R3nF 1 2
Rser 1 3 0.0278586078187
Lser 2 4 3.06758727E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends CSGP_0805_885012007043_3R3nF