.subckt CSGP_0805_885012207014_33nF 1 2
Rser 1 3 0.03079
Lser 2 4 0.00000000030588
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends CSGP_0805_885012207014_33nF