.subckt CSGP_0805_885012207103_1uF 1 2
Rser 1 3 0.0053065272233
Lser 2 4 2.83466289E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends CSGP_0805_885012207103_1uF