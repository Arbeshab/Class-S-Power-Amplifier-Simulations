.subckt CBF_0805_742792036_470ohm 1 2
Rp 1 2 559
Cp 1 2 0.884p
Rs 1 N3 0.3
L1 N3 2 1.4u
.ends CBF_0805_742792036_470ohm