.subckt CSGP_1812_885012010011_4R7nF 1 2
Rser 1 3 0.0944854934425
Lser 2 4 4.17148603E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends CSGP_1812_885012010011_4R7nF
