.subckt 875015119004_150uF 1 2
Rser 1 3 0.00451803569867
Lser 2 4 0.0000000005
C1 3 4 0.00015
Rpar 3 4 66666.6666666667
.ends 875015119004_150uF