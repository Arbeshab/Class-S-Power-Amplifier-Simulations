.subckt CSGP_0805_885012007009_10nF 1 2
Rser 1 3 0.0143302506767
Lser 2 4 2.53788056E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends CSGP_0805_885012007009_10nF