.subckt CSGP_0805_885012007038_0R47nF 1 2
Rser 1 3 0.0888157768288
Lser 2 4 4.59255914E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends CSGP_0805_885012007038_0R47nF