.subckt CSGP_0805_885012007063_1nF 1 2
Rser 1 3 0.0594421507531
Lser 2 4 4.12205624E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends CSGP_0805_885012007063_1nF