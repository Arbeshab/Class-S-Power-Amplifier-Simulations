.subckt CSGP_0805_885012007036_0R22nF 1 2
Rser 1 3 0.115723179071
Lser 2 4 4.36175568E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends CSGP_0805_885012007036_0R22nF