.subckt ASLI_865080545012_100uF 1 2
Rser 1 3 0.31
Lser 2 4 0.000000002805
C1 3 4 0.0001
Rpar 3 4 1000000
.ends ASLI_865080545012_100uF